library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity decodificador is

end entity;

architecture comportamento of decodificador is

begin

end architecture;